module sva_slave(
    input clk,
    input logic rst_n,
    input logic MOSI,
    input logic SS_n,
    input logic tx_valid,
    input logic [7:0] tx_data,
    input logic MISO,
    input logic rx_valid,
    input logic [9:0] rx_data


);
    

endmodule