interface interface_wrapper(clk);
    input clk;
    logic MOSI,MISO,SS_n,rst_n,MISO_ref;
endinterface