package monitor_wrapper;
`include "uvm_macros.svh"
import uvm_pkg::*;
import sequnce_wrapper_item::*;
class monitor_wrapper extends uvm_monitor;
    `uvm_component_utils(monitor_wrapper)
    sequnce_wrapper_item item;
    virtual interface_wrapper if_wrapper;
    uvm_analysis_port #(sequnce_wrapper_item) mon_ap;

    

    function new(string name = "monitor_wrapper", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        // Create the analysis port
        mon_ap = new("mon_ap", this);
    endfunction    

    task run_phase(uvm_phase phase);
        super.run_phase(phase);
        
        forever begin
            item = sequnce_wrapper_item::type_id::create("item");
            // Wait for a valid transaction
           @(negedge if_wrapper.clk);
            
                item.datain = if_wrapper.din;
                item.rx_valid = if_wrapper.rx_valid;
                item.rst_n = if_wrapper.rst_n;
                item.dout = if_wrapper.dout;
                item.tx_valid = if_wrapper.tx_valid;
                
                // Send the item to the analysis export
                mon_ap.write(item);
            end
         
    endtask

endclass //monitor_wrapper extends uvm_monitor;
  
    
endpackage